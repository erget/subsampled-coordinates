netcdf NDVI_example_compacted {
dimensions:
  // NDVI product grid
  lat = 6 ;
  lon = 5 ;
  // Tie points (tp)
  tp_lat = 2 ;
  tp_lon = 2 ;

variables:
  float ndvi(lat, lon) ;
    ndvi : standard_name = "normalized_difference_vegetation_index" ;
    ndvi : interpolation = "tp_interpolation" ;
    ndvi : interpolation_indices = "lat_indices lon_indices" ;
  int lat_indices(tp_lat) ;
    lat_indices : interpolation_dimension = "lat" ;
  int lon_indices(tp_lon) ;
    lon_indices : interpolation_dimension = "lon" ;

  char tp_interpolation ;
    tp_interpolation : interpolation_name = "bi_linear" ;
    tp_interpolation : location_tie_points = "lat lon" ;
  float lat(tp_lat) ;
    lat : standard_name = "latitude" ;
    lat : units = "degrees_north" ;
  float lon(tp_lon) ;
    lon : standard_name = "longitude" ;
    lon : units = "degrees_east" ;

data:
  ndvi =
    0.5119157, 0.04983568, 0.5414233, 0.3076001, 0.8931185,
    0.8581991, 0.7848567, 0.2485297, 0.9762608, 0.4546139,
    0.1063213, 0.8751125, 0.9819403, 0.9346204, 0.2765055,
    0.2011242, 0.7634977, 0.7657007, 0.3465044, 0.9491135,
    0.9431587, 0.04104269, 0.5652257, 0.5340118, 0.8907427,
    0.3514801, 0.1451995, 0.1523716, 0.1563433, 0.7384073 ;
  lat_indices = 0, 5 ;
  lon_indices = 0, 4 ;
  lat = 10, 20 ;
  lon = 10, 30 ;
}
