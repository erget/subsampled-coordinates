��n e t c d f   m w i _ c o m p a c t   {  
 d i m e n s i o n s :  
 	 s c a n l i n e s   =   1 0 0 0   ;  
 	 s c a n p o s       =   1 2 5   ;  
  
 v a r i a b l e s :  
  
                 / /   T w o   b r i g h t n e s s   t e m p e r a t u r e   c h a n n e l s   ( 1 8 . 7   G H z )   u s e   t h e   s a m e   l a t / l o n  
 	 f l o a t   t b 1 8 v ( s c a n l i n e s ,   s c a n p o s )   ;  
 	 	 t b 1 8 v : s t a n d a r d _ n a m e   =   " b r i g h t n e s s _ t e m p e r a t u r e "   ;  
 	 	 t b 1 8 v : t i e _ p o i n t _ i n t e r p o l a t i o n   =   " t i e _ p o i n t s _ 1 8 / i n t e r p o l a t i o n "   ;  
                                 t b 1 8 v : c o o r d i n a t e s   =   " l a t 1 8   l o n 1 8 "  
                 f l o a t   t b 1 8 h ( s c a n l i n e s ,   s c a n p o s )   ;  
 	 	 t b 1 8 h : s t a n d a r d _ n a m e   =   " b r i g h t n e s s _ t e m p e r a t u r e "   ;  
 	 	 t b 1 8 h : t i e _ p o i n t _ i n t e r p o l a t i o n   =   " t i e _ p o i n t s _ 1 8 / i n t e r p o l a t i o n "   ;  
                                 t b 1 8 h : c o o r d i n a t e s   =   " l a t 1 8   l o n 1 8 "  
  
 d a t a :  
  
 g r o u p :   t i e _ p o i n t s _ 1 8   {  
     d i m e n s i o n s :  
     	 s c a n p o s   =   2 5   ;  
     v a r i a b l e s :  
     	 i n t   i n t e r p o l a t i o n   ;  
     	 	 i n t e r p o l a t i o n : t i e _ p o i n t _ i n t e r p o l a t i o n _ n a m e   =   " l i n e a r "   ;  
     	 	 i n t e r p o l a t i o n : t i e _ p o i n t _ i n d i c e s   =   " s c a n p o s _ i n d i c e s "   ;  
     	 	 i n t e r p o l a t i o n : l o c a t i o n _ t i e _ p o i n t s   =   " l a t   l o n "   ;  
     	 i n t   s c a n p o s _ i n d i c e s ( s c a n p o s )   ;  
     	 	 s c a n p o s _ i n d i c e s : l o n g _ n a m e   =   " t i e _ p o i n t _ i n d i c e s _ i n _ i n t e r p o l a t i o n _ d i m e n s i o n "   ;  
     	 	 s c a n p o s _ i n d i c e s : i n t e r p o l a t i o n _ d i m e n s i o n   =   " . . / s c a n p o s "   ;  
     	 f l o a t   l a t 1 8 ( s c a n l i n e s ,   s c a n p o s )   ;  
     	 	 l a t 1 8 : s t a n d a r d _ n a m e   =   " l a t i t u d e "   ;  
     	 	 l a t 1 8 : u n i t s   =   " d e g r e e s _ n o r t h "   ;  
     	 f l o a t   l o n 1 8 ( s c a n l i n e s ,   s c a n p o s )   ;  
     	 	 l o n 1 8 : s t a n d a r d _ n a m e   =   " l o n g i t u d e "   ;  
     	 	 l o n 1 8 : u n i t s   =   " d e g r e e s _ e a s t "   ;  
     d a t a :  
  
       i n t e r p o l a t i o n   =   0   ;  
  
       l a t 1 8   =   f l o a t _ a r r a y ( 1 0 0 0 ,   2 5 )   ;  
  
       l o n 1 8   =   f l o a t _ a r r a y ( 1 0 0 0 ,   2 5 )   ;  
  
       s c a n p o s _ i n d i c e s   =   0 ,   2 4 ,   2 9 ,   . . .   ,   1 2 4  
  
     }   / /   g r o u p   t i e _ p o i n t s  
  
 }  
 