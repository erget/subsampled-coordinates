��n e t c d f   n d v i _ c o m p a c t   {  
 d i m e n s i o n s :  
 	 l a t   =   6   ;  
 	 l o n   =   5   ;  
 v a r i a b l e s :  
 	 f l o a t   n d v i ( l a t ,   l o n )   ;  
 	 	 n d v i : s t a n d a r d _ n a m e   =   " n o r m a l i z e d _ d i f f e r e n c e _ v e g e t a t i o n _ i n d e x "   ;  
 	 	 n d v i : t i e _ p o i n t _ i n t e r p o l a t i o n   =   " t i e _ p o i n t s / i n t e r p o l a t i o n "   ;  
 d a t a :  
  
   n d v i   =  
     0 . 5 1 1 9 1 5 7 ,   0 . 0 4 9 8 3 5 6 8 ,   0 . 5 4 1 4 2 3 3 ,   0 . 3 0 7 6 0 0 1 ,   0 . 8 9 3 1 1 8 5 ,  
     0 . 8 5 8 1 9 9 1 ,   0 . 7 8 4 8 5 6 7 ,   0 . 2 4 8 5 2 9 7 ,   0 . 9 7 6 2 6 0 8 ,   0 . 4 5 4 6 1 3 9 ,  
     0 . 1 0 6 3 2 1 3 ,   0 . 8 7 5 1 1 2 5 ,   0 . 9 8 1 9 4 0 3 ,   0 . 9 3 4 6 2 0 4 ,   0 . 2 7 6 5 0 5 5 ,  
     0 . 2 0 1 1 2 4 2 ,   0 . 7 6 3 4 9 7 7 ,   0 . 7 6 5 7 0 0 7 ,   0 . 3 4 6 5 0 4 4 ,   0 . 9 4 9 1 1 3 5 ,  
     0 . 9 4 3 1 5 8 7 ,   0 . 0 4 1 0 4 2 6 9 ,   0 . 5 6 5 2 2 5 7 ,   0 . 5 3 4 0 1 1 8 ,   0 . 8 9 0 7 4 2 7 ,  
     0 . 3 5 1 4 8 0 1 ,   0 . 1 4 5 1 9 9 5 ,   0 . 1 5 2 3 7 1 6 ,   0 . 1 5 6 3 4 3 3 ,   0 . 7 3 8 4 0 7 3   ;  
  
 g r o u p :   t i e _ p o i n t s   {  
     d i m e n s i o n s :  
     	 l a t   =   2   ;  
     	 l o n   =   2   ;  
     v a r i a b l e s :  
     	 i n t   i n t e r p o l a t i o n   ;  
     	 	 i n t e r p o l a t i o n : t i e _ p o i n t _ i n t e r p o l a t i o n _ n a m e   =   " b i _ l i n e a r "   ;  
     	 	 i n t e r p o l a t i o n : t i e _ p o i n t _ i n d i c e s   =   " l a t _ i n d i c e s   l o n _ i n d i c e s "   ;  
     	 	 i n t e r p o l a t i o n : l o c a t i o n _ t i e _ p o i n t s   =   " l a t   l o n "   ;  
     	 f l o a t   l a t ( l a t )   ;  
     	 	 l a t : s t a n d a r d _ n a m e   =   " l a t i t u d e "   ;  
     	 	 l a t : u n i t s   =   " d e g r e e s _ n o r t h "   ;  
     	 f l o a t   l o n ( l o n )   ;  
     	 	 l o n : s t a n d a r d _ n a m e   =   " l o n g i t u d e "   ;  
     	 	 l o n : u n i t s   =   " d e g r e e s _ e a s t "   ;  
     	 i n t   l a t _ i n d i c e s ( l a t )   ;  
     	 	 l a t _ i n d i c e s : l o n g _ n a m e   =   " t i e _ p o i n t _ i n d i c e s _ i n _ i n t e r p o l a t i o n _ d i m e n s i o n "   ;  
     	 	 l a t _ i n d i c e s : i n t e r p o l a t i o n _ d i m e n s i o n   =   " . . / l a t "   ;  
     	 i n t   l o n _ i n d i c e s ( l o n )   ;  
     	 	 l o n _ i n d i c e s : l o n g _ n a m e   =   " t i e _ p o i n t _ i n d i c e s _ i n _ i n t e r p o l a t i o n _ d i m e n s i o n "   ;  
     	 	 l o n _ i n d i c e s : i n t e r p o l a t i o n _ d i m e n s i o n   =   " . . / l o n "   ;  
     d a t a :  
  
       i n t e r p o l a t i o n   =   0   ;  
  
       l a t   =   1 0 ,   2 0   ;  
  
       l o n   =   1 0 ,   3 0   ;  
  
       l a t _ i n d i c e s   =   0 ,   5   ;  
  
       l o n _ i n d i c e s   =   0 ,   4   ;  
     }   / /   g r o u p   t i e _ p o i n t s  
 }  
 