��n e t c d f   v i i r s _ c o m p a c t   {  
 d i m e n s i o n s :  
 	 t r a c k   =   7 6 8   ;  
 	 s c a n   =   3 2 0 0   ;  
 	 c h a n n e l   =   1 6   ;  
 v a r i a b l e s :  
 	 f l o a t   r a d i a n c e ( t r a c k ,   s c a n ,   c h a n n e l )   ;  
 	 	 r a d i a n c e : t i e _ p o i n t _ i n t e r p o l a t i o n   =   " t p / i n t e r p o l a t i o n "   ;  
 d a t a :  
  
 g r o u p :   t p   {  
     d i m e n s i o n s :  
     	 t r a c k   =   9 6   ;  
     	 s c a n   =   2 0 5   ;  
     	 t r a c k _ i n t e r p o l a t i o n _ z o n e   =   4 8   ;  
     	 s c a n _ i n t e r p o l a t i o n _ z o n e   =   2 0 0   ;  
     v a r i a b l e s :  
     	 i n t   i n t e r p o l a t i o n   ;  
     	 	 i n t e r p o l a t i o n : t i e _ p o i n t _ i n t e r p o l a t i o n _ n a m e   =   " b i _ q u a d r a t i c _ m e t h o d 1 "   ;  
     	 	 i n t e r p o l a t i o n : t i e _ p o i n t _ i n t e r p o l a t i o n _ c o e f f i c i e n t s   =   " e x p a n s i o n _ c o e f f i c i e n t _ t r a c k   a l i g n m e n t _ c o e f f i c i e n t _ t r a c k   e x p a n s i o n _ c o e f f i c i e n t _ s c a n   a l i g n m e n t _ c o e f f i c i e n t _ s c a n "   ;  
     	 	 i n t e r p o l a t i o n : t i e _ p o i n t _ i n t e r p o l a t i o n _ f l a g s   =   " i n t e r p o l a t i o n _ z o n e _ f l a g s "   ;  
     	 	 i n t e r p o l a t i o n : t i e _ p o i n t _ i n d i c e s   =   " t r a c k _ i n d i c e s   s c a n _ i n d i c e s "   ;  
     	 	 i n t e r p o l a t i o n : l o c a t i o n _ t i e _ p o i n t s   =   " l a t   l o n "   ;  
     	 	 i n t e r p o l a t i o n : s e n s o r _ d i r e c t i o n _ t i e _ p o i n t s   =   " s e n _ a z i _ a n g   s e n _ z e n _ a n g "   ;  
     	 	 i n t e r p o l a t i o n : s o l a r _ d i r e c t i o n _ t i e _ p o i n t s   =   " s o l _ a z i _ a n g   s o l _ z e n _ a n g "   ;  
     	 f l o a t   l a t ( t r a c k ,   s c a n )   ;  
     	 	 l a t : s t a n d a r d _ n a m e   =   " l a t i t u d e "   ;  
     	 	 l a t : u n i t s   =   " d e g r e e s _ n o r t h "   ;  
     	 f l o a t   l o n ( t r a c k ,   s c a n )   ;  
     	 	 l o n : s t a n d a r d _ n a m e   =   " l o n g i t u d e "   ;  
     	 	 l o n : u n i t s   =   " d e g r e e s _ e a s t "   ;  
     	 f l o a t   s e n _ a z i _ a n g ( t r a c k ,   s c a n )   ;  
     	 	 s e n _ a z i _ a n g : s t a n d a r d _ n a m e   =   " s e n s o r _ a z i m u t h _ a n g l e "   ;  
     	 	 s e n _ a z i _ a n g : u n i t s   =   " d e g r e e s "   ;  
     	 f l o a t   s e n _ z e n _ a n g ( t r a c k ,   s c a n )   ;  
     	 	 s e n _ z e n _ a n g : s t a n d a r d _ n a m e   =   " s e n s o r _ z e n i t h _ a n g l e "   ;  
     	 	 s e n _ z e n _ a n g : u n i t s   =   " d e g r e e s "   ;  
     	 f l o a t   s o l _ a z i _ a n g ( t r a c k ,   s c a n )   ;  
     	 	 s o l _ a z i _ a n g : s t a n d a r d _ n a m e   =   " s o l a r _ a z i m u t h _ a n g l e "   ;  
     	 	 s o l _ a z i _ a n g : u n i t s   =   " d e g r e e s "   ;  
     	 f l o a t   s o l _ z e n _ a n g ( t r a c k ,   s c a n )   ;  
     	 	 s o l _ z e n _ a n g : s t a n d a r d _ n a m e   =   " s o l a r _ z e n i t h _ a n g l e "   ;  
     	 	 s o l _ z e n _ a n g : u n i t s   =   " d e g r e e s "   ;  
     	 i n t   t r a c k _ i n d i c e s ( t r a c k )   ;  
     	 	 t r a c k _ i n d i c e s : l o n g _ n a m e   =   " t i e _ p o i n t _ i n d i c e s _ i n _ i n t e r p o l a t i o n _ d i m e n s i o n "   ;  
     	 	 t r a c k _ i n d i c e s : i n t e r p o l a t i o n _ d i m e n s i o n   =   " . . / t r a c k "   ;  
     	 i n t   s c a n _ i n d i c e s ( s c a n )   ;  
     	 	 s c a n _ i n d i c e s : l o n g _ n a m e   =   " t i e _ p o i n t _ i n d i c e s _ i n _ i n t e r p o l a t i o n _ d i m e n s i o n "   ;  
     	 	 s c a n _ i n d i c e s : i n t e r p o l a t i o n _ d i m e n s i o n   =   " . . / s c a n "   ;  
     	 s h o r t   e x p a n s i o n _ c o e f f i c i e n t _ t r a c k ( t r a c k _ i n t e r p o l a t i o n _ z o n e ,   s c a n )   ;  
     	 s h o r t   a l i g n m e n t _ c o e f f i c i e n t _ t r a c k ( t r a c k _ i n t e r p o l a t i o n _ z o n e ,   s c a n )   ;  
     	 s h o r t   e x p a n s i o n _ c o e f f i c i e n t _ s c a n ( t r a c k ,   s c a n _ i n t e r p o l a t i o n _ z o n e )   ;  
     	 s h o r t   a l i g n m e n t _ c o e f f i c i e n t _ s c a n ( t r a c k ,   s c a n _ i n t e r p o l a t i o n _ z o n e )   ;  
     	 b y t e   i n t e r p o l a t i o n _ z o n e _ f l a g s ( t r a c k _ i n t e r p o l a t i o n _ z o n e ,   s c a n _ i n t e r p o l a t i o n _ z o n e )   ;  
     	 	 i n t e r p o l a t i o n _ z o n e _ f l a g s : l o n g _ n a m e   =   " i n t e r p o l a t i o n _ c o o r d i n a t e s "   ;  
     	 	 i n t e r p o l a t i o n _ z o n e _ f l a g s : v a l i d _ r a n g e   =   " 1 b ,   7 b "   ;  
     	 	 i n t e r p o l a t i o n _ z o n e _ f l a g s : f l a g _ m a s k s   =   " 1 b ,   2 b ,   4 b "   ;  
     	 	 i n t e r p o l a t i o n _ z o n e _ f l a g s : f l a g _ m e a n i n g s   =   " l o c a t i o n _ u s e _ c a r t e s i a n     s e n s o r _ d i r e c t i o n _ u s e _ c a r t e s i a n     s o l a r _ d i r e c t i o n _ u s e _ c a r t e s i a n "   ;  
     d a t a :  
     }   / /   g r o u p   t p  
 }  
 